entity hello_world is
end hello_world;

architecture one of hello_world is
begin
	process
	begin
		report"Hello world";
	end process;
end one;