entity Transmitter is
  port()